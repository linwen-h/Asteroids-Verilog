module spaceship(clk, reset, start_x, start_y, shooting, direction_x, direction_y, collision, curr_x, curr_y, plot_ship);

input clk, reset, shooting, collision;
input [7:0] start_x;
input [6:0] start_y;

output [7:0] curr_x;
output [6:0] curr_y;



endmodule
