module gameover();
endmodule
