module random_num();
endmodule
