module gameboard();
endmodule
