module main_menu();
endmodule
