module asteroid();

endmodule
